package testing_pkg;
	typedef enum {ADD,SUB,MULT,DIV} opcode_e;
endpackage